`include "16BitAdder.v"

module top;

reg[16:1] a;
reg[16:1] b;
reg cin;
wire[16:1] sum;
wire cout;

	Bit16Adder BA16_0(a, b, cin, sum, cout);

initial
begin
	a[16:1]=16'b0000000000000000;
	#10 b[16:1]=16'b0000000000000000;
	#10 cin=0;
	
	#10 a[16:1]=16'b0000100000100000;b[16:1]=16'b0001000010000011;cin=1;
	#10 a[16:1]=16'b1100000111100000;b[16:1]=16'b0110010000011111;cin=0;
	#10 a[16:1]=16'b0010111100011000;b[16:1]=16'b0011100000110000;cin=0;
	
	#10 a[16:1]=16'b0011110011101110;b[16:1]=16'b0111111111100000;cin=1;
	#10 a[16:1]=16'b0111111100000000;b[16:1]=16'b0000000011110000;cin=0;
	#10 a[16:1]=16'b0111111100000110;b[16:1]=16'b0111000111100000;cin=1;
	
	#10 a[16:1]=16'b1111111111111111;b[16:1]=16'b1111111111111111;cin=1;
	#10;
end

initial
begin
	$monitor($time, ": a = %d, b = %d, cin = %b, Sum = %d, cout = %b", a, b, cin, sum, cout);
	$dumpfile("16BitAdder.vcd");
	$dumpvars;
end

endmodule
